module AHBlite_GPIO_READ( 
    input  wire          HCLK,    
    input  wire          HRESETn, 
    input  wire          HSEL,    
    input  wire   [31:0] HADDR,   
    input  wire    [1:0] HTRANS,  
    input  wire    [2:0] HSIZE,   
    input  wire    [3:0] HPROT,   
    input  wire          HWRITE,  
    input  wire   [31:0] HWDATA,  
    input  wire          HREADY,  
    output wire          HREADYOUT, 
    output wire   [31:0] HRDATA,  
    output wire          HRESP,
    inout  wire   [7:0]  IO_READ
);

assign HRESP = 1'b0;
assign HREADYOUT = 1'b1;

assign HRDATA = {24'b0,IO_READ};
endmodule



